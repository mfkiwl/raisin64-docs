de_isa_def.vh
=============

.. literalinclude:: ../raisin64-cpu/rtl/include/de_isa_def.vh
   :language: verilog
   :linenos:
