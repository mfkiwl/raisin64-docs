io_def.vh
==========

.. literalinclude:: ../raisin64-cpu/rtl/include/io_def.vh
   :language: verilog
   :linenos:
